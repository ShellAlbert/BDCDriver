module led_ctl_by_uart(clk,reset);
endmodule