module rx_fifo(clk,reset,put_pulse,)