module rxclk_sync_to_txclk(clk,reset,)