module pwm_module(clk,reset,pwm1,pwm2);
endmodule
