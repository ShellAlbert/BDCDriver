module rx_bps_module(clk,reset,bps_clk);
endmodule