module rx_module(clk,reset,);
endmodule