module clk_prescale(clk,reset,clk_main);
endmodule