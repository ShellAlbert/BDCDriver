module tb_clk_prescale(clk,clk_out);
endmodule