module H2L_Detect();