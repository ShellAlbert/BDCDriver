module rx_core(clk,reset,H2L_Sig,RXD,);
endmodule